`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // ✅ Bit-level aliases for waveform visibility
  wire t_bit;
  wire q_bit;
  assign t_bit = ui_in[0];
  assign q_bit = uo_out[0];

  // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.vcd");

    // dump everything (keeps your current behavior)
    $dumpvars(0, tb);

    // ✅ force single-bit signals into the VCD so GTKWave can show them
    $dumpvars(1, t_bit);
    $dumpvars(1, q_bit);
    $dumpvars(1, clk);
    $dumpvars(1, rst_n);

    #1;
  end

  // Replace tt_um_example with your module name:
  tt_um_nasser_hadi_tff user_project (

`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
